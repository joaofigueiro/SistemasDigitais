
module BlocoComando(

); 

endmodule; 
