
module BlocoOperativo(

); 

endmodule; 
